`include "baud_gen.sv"
`include "uart_tx.sv"
`include "uart_rx.sv"